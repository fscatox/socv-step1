/**
* Copyright (c) 2023 Politecnico di Torino
*
* This source code is licensed under the BSD-style license found in the
* LICENSE file in the root directory of this source tree.
*
* File              : acc_if.svh
* Author            : Fabio Scatozza <s315216@studenti.polito.it>
* Date              : 13.06.2023
* Last Modified Date: 13.06.2023
* ---------------------------------------------------------------------------
* "acc_if"-related type declarations
*/

`ifndef ACC_IF_SVH
`define ACC_IF_SVH

typedef virtual acc_if.tb v_acctb_if;

`endif

